// look-up table for gf operations
// uses primitive 0x11d, see create_LUT.py
module LUT(index, gf_exp, gf_log);

parameter m = 255;
parameter SIZE = $clog2(m);

input [SIZE-1:0] index;
output [SIZE-1:0] gf_exp, gf_log;

wire [SIZE-1:0] exp_mem[0:255];
wire [SIZE-1:0] log_mem[0:255];

assign gf_exp = exp_mem[index];
assign gf_log = log_mem[index];

assign exp_mem[0] = 1;
assign exp_mem[1] = 2;
assign exp_mem[2] = 4;
assign exp_mem[3] = 8;
assign exp_mem[4] = 16;
assign exp_mem[5] = 32;
assign exp_mem[6] = 64;
assign exp_mem[7] = 128;
assign exp_mem[8] = 29;
assign exp_mem[9] = 58;
assign exp_mem[10] = 116;
assign exp_mem[11] = 232;
assign exp_mem[12] = 205;
assign exp_mem[13] = 135;
assign exp_mem[14] = 19;
assign exp_mem[15] = 38;
assign exp_mem[16] = 76;
assign exp_mem[17] = 152;
assign exp_mem[18] = 45;
assign exp_mem[19] = 90;
assign exp_mem[20] = 180;
assign exp_mem[21] = 117;
assign exp_mem[22] = 234;
assign exp_mem[23] = 201;
assign exp_mem[24] = 143;
assign exp_mem[25] = 3;
assign exp_mem[26] = 6;
assign exp_mem[27] = 12;
assign exp_mem[28] = 24;
assign exp_mem[29] = 48;
assign exp_mem[30] = 96;
assign exp_mem[31] = 192;
assign exp_mem[32] = 157;
assign exp_mem[33] = 39;
assign exp_mem[34] = 78;
assign exp_mem[35] = 156;
assign exp_mem[36] = 37;
assign exp_mem[37] = 74;
assign exp_mem[38] = 148;
assign exp_mem[39] = 53;
assign exp_mem[40] = 106;
assign exp_mem[41] = 212;
assign exp_mem[42] = 181;
assign exp_mem[43] = 119;
assign exp_mem[44] = 238;
assign exp_mem[45] = 193;
assign exp_mem[46] = 159;
assign exp_mem[47] = 35;
assign exp_mem[48] = 70;
assign exp_mem[49] = 140;
assign exp_mem[50] = 5;
assign exp_mem[51] = 10;
assign exp_mem[52] = 20;
assign exp_mem[53] = 40;
assign exp_mem[54] = 80;
assign exp_mem[55] = 160;
assign exp_mem[56] = 93;
assign exp_mem[57] = 186;
assign exp_mem[58] = 105;
assign exp_mem[59] = 210;
assign exp_mem[60] = 185;
assign exp_mem[61] = 111;
assign exp_mem[62] = 222;
assign exp_mem[63] = 161;
assign exp_mem[64] = 95;
assign exp_mem[65] = 190;
assign exp_mem[66] = 97;
assign exp_mem[67] = 194;
assign exp_mem[68] = 153;
assign exp_mem[69] = 47;
assign exp_mem[70] = 94;
assign exp_mem[71] = 188;
assign exp_mem[72] = 101;
assign exp_mem[73] = 202;
assign exp_mem[74] = 137;
assign exp_mem[75] = 15;
assign exp_mem[76] = 30;
assign exp_mem[77] = 60;
assign exp_mem[78] = 120;
assign exp_mem[79] = 240;
assign exp_mem[80] = 253;
assign exp_mem[81] = 231;
assign exp_mem[82] = 211;
assign exp_mem[83] = 187;
assign exp_mem[84] = 107;
assign exp_mem[85] = 214;
assign exp_mem[86] = 177;
assign exp_mem[87] = 127;
assign exp_mem[88] = 254;
assign exp_mem[89] = 225;
assign exp_mem[90] = 223;
assign exp_mem[91] = 163;
assign exp_mem[92] = 91;
assign exp_mem[93] = 182;
assign exp_mem[94] = 113;
assign exp_mem[95] = 226;
assign exp_mem[96] = 217;
assign exp_mem[97] = 175;
assign exp_mem[98] = 67;
assign exp_mem[99] = 134;
assign exp_mem[100] = 17;
assign exp_mem[101] = 34;
assign exp_mem[102] = 68;
assign exp_mem[103] = 136;
assign exp_mem[104] = 13;
assign exp_mem[105] = 26;
assign exp_mem[106] = 52;
assign exp_mem[107] = 104;
assign exp_mem[108] = 208;
assign exp_mem[109] = 189;
assign exp_mem[110] = 103;
assign exp_mem[111] = 206;
assign exp_mem[112] = 129;
assign exp_mem[113] = 31;
assign exp_mem[114] = 62;
assign exp_mem[115] = 124;
assign exp_mem[116] = 248;
assign exp_mem[117] = 237;
assign exp_mem[118] = 199;
assign exp_mem[119] = 147;
assign exp_mem[120] = 59;
assign exp_mem[121] = 118;
assign exp_mem[122] = 236;
assign exp_mem[123] = 197;
assign exp_mem[124] = 151;
assign exp_mem[125] = 51;
assign exp_mem[126] = 102;
assign exp_mem[127] = 204;
assign exp_mem[128] = 133;
assign exp_mem[129] = 23;
assign exp_mem[130] = 46;
assign exp_mem[131] = 92;
assign exp_mem[132] = 184;
assign exp_mem[133] = 109;
assign exp_mem[134] = 218;
assign exp_mem[135] = 169;
assign exp_mem[136] = 79;
assign exp_mem[137] = 158;
assign exp_mem[138] = 33;
assign exp_mem[139] = 66;
assign exp_mem[140] = 132;
assign exp_mem[141] = 21;
assign exp_mem[142] = 42;
assign exp_mem[143] = 84;
assign exp_mem[144] = 168;
assign exp_mem[145] = 77;
assign exp_mem[146] = 154;
assign exp_mem[147] = 41;
assign exp_mem[148] = 82;
assign exp_mem[149] = 164;
assign exp_mem[150] = 85;
assign exp_mem[151] = 170;
assign exp_mem[152] = 73;
assign exp_mem[153] = 146;
assign exp_mem[154] = 57;
assign exp_mem[155] = 114;
assign exp_mem[156] = 228;
assign exp_mem[157] = 213;
assign exp_mem[158] = 183;
assign exp_mem[159] = 115;
assign exp_mem[160] = 230;
assign exp_mem[161] = 209;
assign exp_mem[162] = 191;
assign exp_mem[163] = 99;
assign exp_mem[164] = 198;
assign exp_mem[165] = 145;
assign exp_mem[166] = 63;
assign exp_mem[167] = 126;
assign exp_mem[168] = 252;
assign exp_mem[169] = 229;
assign exp_mem[170] = 215;
assign exp_mem[171] = 179;
assign exp_mem[172] = 123;
assign exp_mem[173] = 246;
assign exp_mem[174] = 241;
assign exp_mem[175] = 255;
assign exp_mem[176] = 227;
assign exp_mem[177] = 219;
assign exp_mem[178] = 171;
assign exp_mem[179] = 75;
assign exp_mem[180] = 150;
assign exp_mem[181] = 49;
assign exp_mem[182] = 98;
assign exp_mem[183] = 196;
assign exp_mem[184] = 149;
assign exp_mem[185] = 55;
assign exp_mem[186] = 110;
assign exp_mem[187] = 220;
assign exp_mem[188] = 165;
assign exp_mem[189] = 87;
assign exp_mem[190] = 174;
assign exp_mem[191] = 65;
assign exp_mem[192] = 130;
assign exp_mem[193] = 25;
assign exp_mem[194] = 50;
assign exp_mem[195] = 100;
assign exp_mem[196] = 200;
assign exp_mem[197] = 141;
assign exp_mem[198] = 7;
assign exp_mem[199] = 14;
assign exp_mem[200] = 28;
assign exp_mem[201] = 56;
assign exp_mem[202] = 112;
assign exp_mem[203] = 224;
assign exp_mem[204] = 221;
assign exp_mem[205] = 167;
assign exp_mem[206] = 83;
assign exp_mem[207] = 166;
assign exp_mem[208] = 81;
assign exp_mem[209] = 162;
assign exp_mem[210] = 89;
assign exp_mem[211] = 178;
assign exp_mem[212] = 121;
assign exp_mem[213] = 242;
assign exp_mem[214] = 249;
assign exp_mem[215] = 239;
assign exp_mem[216] = 195;
assign exp_mem[217] = 155;
assign exp_mem[218] = 43;
assign exp_mem[219] = 86;
assign exp_mem[220] = 172;
assign exp_mem[221] = 69;
assign exp_mem[222] = 138;
assign exp_mem[223] = 9;
assign exp_mem[224] = 18;
assign exp_mem[225] = 36;
assign exp_mem[226] = 72;
assign exp_mem[227] = 144;
assign exp_mem[228] = 61;
assign exp_mem[229] = 122;
assign exp_mem[230] = 244;
assign exp_mem[231] = 245;
assign exp_mem[232] = 247;
assign exp_mem[233] = 243;
assign exp_mem[234] = 251;
assign exp_mem[235] = 235;
assign exp_mem[236] = 203;
assign exp_mem[237] = 139;
assign exp_mem[238] = 11;
assign exp_mem[239] = 22;
assign exp_mem[240] = 44;
assign exp_mem[241] = 88;
assign exp_mem[242] = 176;
assign exp_mem[243] = 125;
assign exp_mem[244] = 250;
assign exp_mem[245] = 233;
assign exp_mem[246] = 207;
assign exp_mem[247] = 131;
assign exp_mem[248] = 27;
assign exp_mem[249] = 54;
assign exp_mem[250] = 108;
assign exp_mem[251] = 216;
assign exp_mem[252] = 173;
assign exp_mem[253] = 71;
assign exp_mem[254] = 142;
assign exp_mem[255] = 1;

assign log_mem[0] = 0;
assign log_mem[1] = 0;
assign log_mem[2] = 1;
assign log_mem[3] = 25;
assign log_mem[4] = 2;
assign log_mem[5] = 50;
assign log_mem[6] = 26;
assign log_mem[7] = 198;
assign log_mem[8] = 3;
assign log_mem[9] = 223;
assign log_mem[10] = 51;
assign log_mem[11] = 238;
assign log_mem[12] = 27;
assign log_mem[13] = 104;
assign log_mem[14] = 199;
assign log_mem[15] = 75;
assign log_mem[16] = 4;
assign log_mem[17] = 100;
assign log_mem[18] = 224;
assign log_mem[19] = 14;
assign log_mem[20] = 52;
assign log_mem[21] = 141;
assign log_mem[22] = 239;
assign log_mem[23] = 129;
assign log_mem[24] = 28;
assign log_mem[25] = 193;
assign log_mem[26] = 105;
assign log_mem[27] = 248;
assign log_mem[28] = 200;
assign log_mem[29] = 8;
assign log_mem[30] = 76;
assign log_mem[31] = 113;
assign log_mem[32] = 5;
assign log_mem[33] = 138;
assign log_mem[34] = 101;
assign log_mem[35] = 47;
assign log_mem[36] = 225;
assign log_mem[37] = 36;
assign log_mem[38] = 15;
assign log_mem[39] = 33;
assign log_mem[40] = 53;
assign log_mem[41] = 147;
assign log_mem[42] = 142;
assign log_mem[43] = 218;
assign log_mem[44] = 240;
assign log_mem[45] = 18;
assign log_mem[46] = 130;
assign log_mem[47] = 69;
assign log_mem[48] = 29;
assign log_mem[49] = 181;
assign log_mem[50] = 194;
assign log_mem[51] = 125;
assign log_mem[52] = 106;
assign log_mem[53] = 39;
assign log_mem[54] = 249;
assign log_mem[55] = 185;
assign log_mem[56] = 201;
assign log_mem[57] = 154;
assign log_mem[58] = 9;
assign log_mem[59] = 120;
assign log_mem[60] = 77;
assign log_mem[61] = 228;
assign log_mem[62] = 114;
assign log_mem[63] = 166;
assign log_mem[64] = 6;
assign log_mem[65] = 191;
assign log_mem[66] = 139;
assign log_mem[67] = 98;
assign log_mem[68] = 102;
assign log_mem[69] = 221;
assign log_mem[70] = 48;
assign log_mem[71] = 253;
assign log_mem[72] = 226;
assign log_mem[73] = 152;
assign log_mem[74] = 37;
assign log_mem[75] = 179;
assign log_mem[76] = 16;
assign log_mem[77] = 145;
assign log_mem[78] = 34;
assign log_mem[79] = 136;
assign log_mem[80] = 54;
assign log_mem[81] = 208;
assign log_mem[82] = 148;
assign log_mem[83] = 206;
assign log_mem[84] = 143;
assign log_mem[85] = 150;
assign log_mem[86] = 219;
assign log_mem[87] = 189;
assign log_mem[88] = 241;
assign log_mem[89] = 210;
assign log_mem[90] = 19;
assign log_mem[91] = 92;
assign log_mem[92] = 131;
assign log_mem[93] = 56;
assign log_mem[94] = 70;
assign log_mem[95] = 64;
assign log_mem[96] = 30;
assign log_mem[97] = 66;
assign log_mem[98] = 182;
assign log_mem[99] = 163;
assign log_mem[100] = 195;
assign log_mem[101] = 72;
assign log_mem[102] = 126;
assign log_mem[103] = 110;
assign log_mem[104] = 107;
assign log_mem[105] = 58;
assign log_mem[106] = 40;
assign log_mem[107] = 84;
assign log_mem[108] = 250;
assign log_mem[109] = 133;
assign log_mem[110] = 186;
assign log_mem[111] = 61;
assign log_mem[112] = 202;
assign log_mem[113] = 94;
assign log_mem[114] = 155;
assign log_mem[115] = 159;
assign log_mem[116] = 10;
assign log_mem[117] = 21;
assign log_mem[118] = 121;
assign log_mem[119] = 43;
assign log_mem[120] = 78;
assign log_mem[121] = 212;
assign log_mem[122] = 229;
assign log_mem[123] = 172;
assign log_mem[124] = 115;
assign log_mem[125] = 243;
assign log_mem[126] = 167;
assign log_mem[127] = 87;
assign log_mem[128] = 7;
assign log_mem[129] = 112;
assign log_mem[130] = 192;
assign log_mem[131] = 247;
assign log_mem[132] = 140;
assign log_mem[133] = 128;
assign log_mem[134] = 99;
assign log_mem[135] = 13;
assign log_mem[136] = 103;
assign log_mem[137] = 74;
assign log_mem[138] = 222;
assign log_mem[139] = 237;
assign log_mem[140] = 49;
assign log_mem[141] = 197;
assign log_mem[142] = 254;
assign log_mem[143] = 24;
assign log_mem[144] = 227;
assign log_mem[145] = 165;
assign log_mem[146] = 153;
assign log_mem[147] = 119;
assign log_mem[148] = 38;
assign log_mem[149] = 184;
assign log_mem[150] = 180;
assign log_mem[151] = 124;
assign log_mem[152] = 17;
assign log_mem[153] = 68;
assign log_mem[154] = 146;
assign log_mem[155] = 217;
assign log_mem[156] = 35;
assign log_mem[157] = 32;
assign log_mem[158] = 137;
assign log_mem[159] = 46;
assign log_mem[160] = 55;
assign log_mem[161] = 63;
assign log_mem[162] = 209;
assign log_mem[163] = 91;
assign log_mem[164] = 149;
assign log_mem[165] = 188;
assign log_mem[166] = 207;
assign log_mem[167] = 205;
assign log_mem[168] = 144;
assign log_mem[169] = 135;
assign log_mem[170] = 151;
assign log_mem[171] = 178;
assign log_mem[172] = 220;
assign log_mem[173] = 252;
assign log_mem[174] = 190;
assign log_mem[175] = 97;
assign log_mem[176] = 242;
assign log_mem[177] = 86;
assign log_mem[178] = 211;
assign log_mem[179] = 171;
assign log_mem[180] = 20;
assign log_mem[181] = 42;
assign log_mem[182] = 93;
assign log_mem[183] = 158;
assign log_mem[184] = 132;
assign log_mem[185] = 60;
assign log_mem[186] = 57;
assign log_mem[187] = 83;
assign log_mem[188] = 71;
assign log_mem[189] = 109;
assign log_mem[190] = 65;
assign log_mem[191] = 162;
assign log_mem[192] = 31;
assign log_mem[193] = 45;
assign log_mem[194] = 67;
assign log_mem[195] = 216;
assign log_mem[196] = 183;
assign log_mem[197] = 123;
assign log_mem[198] = 164;
assign log_mem[199] = 118;
assign log_mem[200] = 196;
assign log_mem[201] = 23;
assign log_mem[202] = 73;
assign log_mem[203] = 236;
assign log_mem[204] = 127;
assign log_mem[205] = 12;
assign log_mem[206] = 111;
assign log_mem[207] = 246;
assign log_mem[208] = 108;
assign log_mem[209] = 161;
assign log_mem[210] = 59;
assign log_mem[211] = 82;
assign log_mem[212] = 41;
assign log_mem[213] = 157;
assign log_mem[214] = 85;
assign log_mem[215] = 170;
assign log_mem[216] = 251;
assign log_mem[217] = 96;
assign log_mem[218] = 134;
assign log_mem[219] = 177;
assign log_mem[220] = 187;
assign log_mem[221] = 204;
assign log_mem[222] = 62;
assign log_mem[223] = 90;
assign log_mem[224] = 203;
assign log_mem[225] = 89;
assign log_mem[226] = 95;
assign log_mem[227] = 176;
assign log_mem[228] = 156;
assign log_mem[229] = 169;
assign log_mem[230] = 160;
assign log_mem[231] = 81;
assign log_mem[232] = 11;
assign log_mem[233] = 245;
assign log_mem[234] = 22;
assign log_mem[235] = 235;
assign log_mem[236] = 122;
assign log_mem[237] = 117;
assign log_mem[238] = 44;
assign log_mem[239] = 215;
assign log_mem[240] = 79;
assign log_mem[241] = 174;
assign log_mem[242] = 213;
assign log_mem[243] = 233;
assign log_mem[244] = 230;
assign log_mem[245] = 231;
assign log_mem[246] = 173;
assign log_mem[247] = 232;
assign log_mem[248] = 116;
assign log_mem[249] = 214;
assign log_mem[250] = 244;
assign log_mem[251] = 234;
assign log_mem[252] = 168;
assign log_mem[253] = 80;
assign log_mem[254] = 88;
assign log_mem[255] = 175;

endmodule
