module my_dff;
